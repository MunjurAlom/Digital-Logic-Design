CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 60 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 237 271 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9281 0 0
2
43727 0
0
13 Logic Switch~
5 239 218 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8464 0 0
2
43727 0
0
13 Logic Switch~
5 236 168 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7168 0 0
2
43727 0
0
9 Inverter~
13 349 281 0 2 22
0 3 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3171 0 0
2
43727 0
0
8 4-In OR~
219 801 532 0 5 22
0 8 7 6 5 4
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U4B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
4139 0 0
2
43727 0
0
5 7415~
219 607 637 0 4 22
0 10 9 3 5
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 5 0
1 U
6435 0 0
2
43727 0
0
5 7415~
219 604 580 0 4 22
0 10 9 2 6
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 5 0
1 U
5283 0 0
2
43727 0
0
5 7415~
219 604 521 0 4 22
0 10 11 3 7
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 3 0
1 U
6874 0 0
2
43727 0
0
5 7415~
219 604 465 0 4 22
0 12 9 3 8
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
5305 0 0
2
43727 0
0
14 Logic Display~
6 980 490 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
34 0 0
2
43727 0
0
14 Logic Display~
6 901 243 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
969 0 0
2
43727 0
0
8 4-In OR~
219 790 272 0 5 22
0 17 16 15 14 13
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
8402 0 0
2
43727 0
0
5 7415~
219 601 379 0 4 22
0 10 9 3 14
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
3751 0 0
2
43727 0
0
5 7415~
219 599 311 0 4 22
0 10 11 2 15
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 2 0
1 U
4292 0 0
2
43727 0
0
5 7415~
219 596 250 0 4 22
0 12 9 2 16
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 2 0
1 U
6118 0 0
2
43727 0
0
5 7415~
219 595 183 0 4 22
0 12 11 3 17
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 2 0
1 U
34 0 0
2
43727 0
0
9 Inverter~
13 360 218 0 2 22
0 9 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
6357 0 0
2
43727 0
0
9 Inverter~
13 360 168 0 2 22
0 10 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
319 0 0
2
43727 0
0
37
3 0 2 0 0 8320 0 7 0 0 3 3
580 589
438 589
438 281
0 3 2 0 0 0 0 0 14 3 0 3
530 281
530 320
575 320
2 3 2 0 0 0 0 4 15 0 0 4
370 281
564 281
564 259
572 259
0 3 3 0 0 8192 0 0 16 5 0 4
326 271
326 235
571 235
571 192
1 1 3 0 0 0 0 1 4 0 0 4
249 271
326 271
326 281
334 281
5 1 4 0 0 4224 0 5 10 0 0 3
834 532
980 532
980 508
4 4 5 0 0 4224 0 6 5 0 0 4
628 637
771 637
771 546
784 546
4 3 6 0 0 4224 0 7 5 0 0 4
625 580
752 580
752 537
784 537
4 2 7 0 0 4224 0 8 5 0 0 4
625 521
776 521
776 528
784 528
4 1 8 0 0 4224 0 9 5 0 0 4
625 465
776 465
776 519
784 519
0 3 3 0 0 0 0 0 6 19 0 3
430 474
430 646
583 646
0 2 9 0 0 4096 0 0 6 20 0 3
467 465
467 637
583 637
0 1 10 0 0 4096 0 0 6 18 0 3
483 512
483 628
583 628
0 2 9 0 0 0 0 0 7 20 0 3
502 465
502 580
580 580
0 1 10 0 0 0 0 0 7 18 0 3
526 512
526 571
580 571
0 3 3 0 0 0 0 0 8 19 0 3
538 474
538 530
580 530
0 2 11 0 0 4224 0 0 8 30 0 3
551 311
551 521
580 521
0 1 10 0 0 8192 0 0 8 27 0 3
386 370
386 512
580 512
0 3 3 0 0 0 0 0 9 28 0 3
411 388
411 474
580 474
0 2 9 0 0 0 0 0 9 29 0 3
434 379
434 465
580 465
0 1 12 0 0 4224 0 0 9 35 0 3
458 170
458 456
580 456
5 1 13 0 0 4224 0 12 11 0 0 3
823 272
901 272
901 261
4 4 14 0 0 4224 0 13 12 0 0 4
622 379
760 379
760 286
773 286
4 3 15 0 0 4224 0 14 12 0 0 4
620 311
733 311
733 277
773 277
4 2 16 0 0 4224 0 15 12 0 0 4
617 250
760 250
760 268
773 268
4 1 17 0 0 4224 0 16 12 0 0 4
616 183
765 183
765 259
773 259
0 1 10 0 0 8320 0 0 13 37 0 3
302 168
302 370
577 370
0 3 3 0 0 8320 0 0 13 5 0 3
264 271
264 388
577 388
0 2 9 0 0 8320 0 0 13 36 0 3
291 218
291 379
577 379
0 2 11 0 0 0 0 0 14 34 0 3
497 183
497 311
575 311
0 1 10 0 0 0 0 0 14 37 0 3
322 168
322 302
575 302
0 2 9 0 0 0 0 0 15 36 0 3
341 218
341 250
572 250
0 1 12 0 0 0 0 0 15 35 0 3
531 170
531 241
572 241
2 2 11 0 0 0 0 17 16 0 0 3
381 218
381 183
571 183
2 1 12 0 0 0 0 18 16 0 0 4
381 168
381 170
571 170
571 174
1 1 9 0 0 0 0 2 17 0 0 2
251 218
345 218
1 1 10 0 0 0 0 3 18 0 0 2
248 168
345 168
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
878 498 939 522
888 506 928 522
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
835 241 880 265
845 249 869 265
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
412 93 577 117
422 101 566 117
18 Full Adder Circuit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
176 260 205 284
186 268 194 284
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
174 201 203 225
184 209 192 225
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
171 149 200 173
181 157 189 173
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
