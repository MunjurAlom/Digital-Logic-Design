CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 192 358 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43727.5 0
0
13 Logic Switch~
5 199 200 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43727.5 0
0
13 Logic Switch~
5 199 264 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
43727.5 0
0
13 Logic Switch~
5 196 148 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
43727.5 0
0
14 Logic Display~
6 843 134 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
43727.5 0
0
9 2-In NOR~
219 559 246 0 3 22
0 2 6 3
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5572 0 0
2
43727.5 0
0
9 2-In NOR~
219 552 166 0 3 22
0 7 3 4
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8901 0 0
2
43727.5 0
0
9 2-In AND~
219 352 255 0 3 22
0 5 8 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7361 0 0
2
43727.5 0
0
9 2-In AND~
219 346 157 0 3 22
0 9 5 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4747 0 0
2
43727.5 0
0
9
1 1 2 0 0 12432 0 6 1 0 0 4
546 237
440 237
440 358
204 358
3 2 3 0 0 12416 0 6 7 0 0 6
598 246
602 246
602 186
531 186
531 175
539 175
3 1 4 0 0 4224 0 7 5 0 0 3
591 166
843 166
843 152
1 0 5 0 0 4096 0 2 0 0 9 2
211 200
288 200
3 2 6 0 0 4224 0 8 6 0 0 2
373 255
546 255
3 1 7 0 0 4224 0 9 7 0 0 2
367 157
539 157
1 2 8 0 0 4224 0 3 8 0 0 2
211 264
328 264
1 1 9 0 0 4224 0 4 9 0 0 2
208 148
322 148
1 2 5 0 0 8320 0 8 9 0 0 4
328 246
288 246
288 166
322 166
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
340 77 457 101
350 85 446 101
12 SR Flip Flop
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
136 347 165 371
146 355 154 371
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
139 187 176 211
149 195 165 211
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
132 248 161 272
142 256 150 272
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
130 132 159 156
140 140 148 156
1 R
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
