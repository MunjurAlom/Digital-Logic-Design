CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 195 253 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3472 0 0
2
43726.9 0
0
13 Logic Switch~
5 196 170 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9998 0 0
2
43726.9 0
0
14 Logic Display~
6 679 392 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
43726.9 0
0
9 2-In AND~
219 509 405 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4597 0 0
2
43726.9 0
0
14 Logic Display~
6 826 171 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
43726.9 0
0
8 2-In OR~
219 621 201 0 3 22
0 7 6 5
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3670 0 0
2
43726.9 0
0
9 2-In AND~
219 466 273 0 3 22
0 4 8 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5616 0 0
2
43726.9 0
0
9 2-In AND~
219 465 167 0 3 22
0 9 3 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9323 0 0
2
43726.9 0
0
9 Inverter~
13 334 253 0 2 22
0 3 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
317 0 0
2
43726.9 0
0
9 Inverter~
13 333 167 0 2 22
0 4 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3108 0 0
2
43726.9 0
0
12
3 1 2 0 0 4224 0 4 3 0 0 5
530 405
667 405
667 418
679 418
679 410
0 2 3 0 0 8320 0 0 4 11 0 3
250 253
250 414
485 414
0 1 4 0 0 4096 0 0 4 8 0 3
404 268
404 396
485 396
3 1 5 0 0 4224 0 6 5 0 0 5
654 201
782 201
782 208
826 208
826 189
3 2 6 0 0 4224 0 7 6 0 0 4
487 273
600 273
600 210
608 210
3 1 7 0 0 4224 0 8 6 0 0 4
486 167
600 167
600 192
608 192
2 2 8 0 0 4224 0 9 7 0 0 4
355 253
429 253
429 282
442 282
0 1 4 0 0 8320 0 0 7 12 0 5
277 170
277 268
434 268
434 264
442 264
0 2 3 0 0 0 0 0 8 11 0 5
305 253
305 182
433 182
433 176
441 176
2 1 9 0 0 4224 0 10 8 0 0 4
354 167
433 167
433 158
441 158
1 1 3 0 0 0 0 1 9 0 0 2
207 253
319 253
1 1 4 0 0 0 0 2 10 0 0 4
208 170
310 170
310 167
318 167
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
318 32 483 56
328 40 472 56
18 Half Adder Circuit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
701 164 746 188
711 172 735 188
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
556 370 625 394
566 378 614 394
6 Carray
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
485 238 530 262
495 246 519 262
3 AB'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
480 114 525 138
490 122 514 138
3 A'B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
355 229 392 253
365 237 381 253
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
364 145 401 169
374 153 390 169
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
146 235 175 259
156 243 164 259
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
146 150 175 174
156 158 164 174
1 A
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
