CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 156 342 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43727.9 0
0
13 Logic Switch~
5 167 258 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89908e-315 0
0
13 Logic Switch~
5 165 208 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89908e-315 5.26354e-315
0
13 Logic Switch~
5 165 151 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89908e-315 5.30499e-315
0
14 Logic Display~
6 718 131 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89908e-315 5.32571e-315
0
9 2-In NOR~
219 549 248 0 3 22
0 2 8 3
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5572 0 0
2
5.89908e-315 5.34643e-315
0
9 2-In NOR~
219 548 153 0 3 22
0 9 3 4
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8901 0 0
2
5.89908e-315 5.3568e-315
0
5 7415~
219 364 257 0 4 22
0 5 6 3 8
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
7361 0 0
2
5.89908e-315 5.36716e-315
0
5 7415~
219 358 150 0 4 22
0 4 7 5 9
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
4747 0 0
2
5.89908e-315 5.37752e-315
0
11
1 1 2 0 0 4224 0 1 6 0 0 4
168 342
528 342
528 239
536 239
3 0 3 0 0 12416 0 8 0 0 5 5
340 266
336 266
336 303
627 303
627 248
1 0 4 0 0 12416 0 9 0 0 4 5
334 141
330 141
330 114
611 114
611 153
3 1 4 0 0 0 0 7 5 0 0 3
587 153
718 153
718 149
2 3 3 0 0 0 0 7 6 0 0 6
535 162
522 162
522 210
680 210
680 248
588 248
1 0 5 0 0 4224 0 3 0 0 7 2
177 208
301 208
3 1 5 0 0 0 0 9 8 0 0 4
334 159
301 159
301 248
340 248
1 2 6 0 0 8320 0 2 8 0 0 3
179 258
179 257
340 257
1 2 7 0 0 8320 0 4 9 0 0 3
177 151
177 150
334 150
4 2 8 0 0 4224 0 8 6 0 0 2
385 257
536 257
4 1 9 0 0 4224 0 9 7 0 0 4
379 150
527 150
527 144
535 144
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
314 33 431 57
324 41 420 57
12 JK Flip Flop
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
106 135 135 159
116 143 124 159
1 k
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
100 186 137 210
110 194 126 210
2 cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
106 240 135 264
116 248 124 264
1 j
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
