CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 122 192 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
317 0 0
2
43728 0
0
13 Logic Switch~
5 120 145 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3108 0 0
2
43728 0
0
13 Logic Switch~
5 117 96 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4299 0 0
2
43728 0
0
9 Inverter~
13 227 192 0 2 22
0 7 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
9672 0 0
2
43728 0
0
9 Inverter~
13 226 145 0 2 22
0 8 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
7876 0 0
2
43728 0
0
9 Inverter~
13 226 96 0 2 22
0 9 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
6369 0 0
2
43728 0
0
8 4-In OR~
219 615 379 0 5 22
0 6 5 4 3 2
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U4B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
9172 0 0
2
43728 0
0
8 4-In OR~
219 554 148 0 5 22
0 17 16 15 14 13
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
7100 0 0
2
43728 0
0
14 Logic Display~
6 750 334 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3820 0 0
2
43728 0
0
5 7415~
219 444 447 0 4 22
0 9 8 7 3
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
7678 0 0
2
43728 0
0
5 7415~
219 443 404 0 4 22
0 9 11 10 4
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
961 0 0
2
43728 0
0
5 7415~
219 443 361 0 4 22
0 12 8 10 5
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 2 0
1 U
3178 0 0
2
43728 0
0
5 7415~
219 441 321 0 4 22
0 12 11 7 6
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 2 0
1 U
3409 0 0
2
43728 0
0
5 7415~
219 441 240 0 4 22
0 9 8 7 14
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 2 0
1 U
3951 0 0
2
43728 0
0
5 7415~
219 441 194 0 4 22
0 12 8 7 15
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 1 0
1 U
8885 0 0
2
43728 0
0
5 7415~
219 440 148 0 4 22
0 12 8 10 16
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
3780 0 0
2
43728 0
0
5 7415~
219 440 106 0 4 22
0 12 11 7 17
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
9265 0 0
2
43728 0
0
14 Logic Display~
6 758 106 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9442 0 0
2
43728 0
0
37
5 1 2 0 0 4224 0 7 9 0 0 3
648 379
750 379
750 352
4 4 3 0 0 12432 0 7 10 0 0 4
598 393
594 393
594 447
465 447
4 3 4 0 0 4224 0 11 7 0 0 4
464 404
590 404
590 384
598 384
4 2 5 0 0 4224 0 12 7 0 0 4
464 361
585 361
585 375
598 375
4 1 6 0 0 4224 0 13 7 0 0 4
462 321
590 321
590 366
598 366
0 3 7 0 0 8192 0 0 10 23 0 3
196 249
196 456
420 456
0 2 8 0 0 4096 0 0 10 24 0 3
214 240
214 447
420 447
0 1 9 0 0 4096 0 0 10 25 0 3
239 231
239 438
420 438
0 3 10 0 0 8192 0 0 11 12 0 3
343 370
343 413
419 413
0 2 11 0 0 4096 0 0 11 16 0 3
351 321
351 404
419 404
0 1 9 0 0 0 0 0 11 25 0 3
357 231
357 395
419 395
0 3 10 0 0 4224 0 0 12 29 0 3
258 192
258 370
419 370
0 2 8 0 0 0 0 0 12 24 0 3
375 240
375 361
419 361
0 1 12 0 0 4096 0 0 12 17 0 3
388 312
388 352
419 352
0 3 7 0 0 0 0 0 13 23 0 3
280 249
280 330
417 330
0 2 11 0 0 4224 0 0 13 33 0 3
290 145
290 321
417 321
0 1 12 0 0 4224 0 0 13 34 0 3
312 96
312 312
417 312
5 1 13 0 0 4224 0 8 18 0 0 3
587 148
758 148
758 124
4 4 14 0 0 8320 0 14 8 0 0 4
462 240
524 240
524 162
537 162
4 3 15 0 0 4224 0 15 8 0 0 4
462 194
513 194
513 153
537 153
4 2 16 0 0 4224 0 16 8 0 0 4
461 148
529 148
529 144
537 144
4 1 17 0 0 4224 0 17 8 0 0 4
461 106
529 106
529 135
537 135
0 3 7 0 0 8320 0 0 14 35 0 3
165 192
165 249
417 249
0 2 8 0 0 8320 0 0 14 36 0 3
180 145
180 240
417 240
0 1 9 0 0 8320 0 0 14 37 0 3
198 96
198 231
417 231
0 3 7 0 0 0 0 0 15 35 0 5
192 192
192 210
409 210
409 203
417 203
0 2 8 0 0 0 0 0 15 30 0 4
326 160
326 197
417 197
417 194
0 1 12 0 0 0 0 0 15 34 0 3
350 96
350 185
417 185
2 3 10 0 0 0 0 4 16 0 0 4
248 192
403 192
403 157
416 157
0 2 8 0 0 0 0 0 16 36 0 5
205 145
205 160
338 160
338 148
416 148
0 1 12 0 0 0 0 0 16 34 0 3
384 96
384 139
416 139
0 3 7 0 0 0 0 0 17 35 0 5
203 192
203 170
303 170
303 115
416 115
2 2 11 0 0 0 0 5 17 0 0 4
247 145
293 145
293 106
416 106
2 1 12 0 0 0 0 6 17 0 0 4
247 96
408 96
408 97
416 97
1 1 7 0 0 0 0 1 4 0 0 2
134 192
212 192
1 1 8 0 0 0 0 2 5 0 0 2
132 145
211 145
1 1 9 0 0 0 0 3 6 0 0 2
129 96
211 96
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
312 19 461 43
322 27 450 43
16 Full Subtraction
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
629 115 682 139
639 123 671 139
4 Brow
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
667 347 712 371
677 355 701 371
3 SUB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
77 177 106 201
87 185 95 201
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
82 129 111 153
92 137 100 153
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
74 76 103 100
84 84 92 100
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
